
`timescale 1 ns / 1 ps
    module p_ram_t # (
        parameter DATA_WIDTH = 3,
        parameter ADDR_WIDTH = 10
    ) (
        input wire clk,
        input wire [ADDR_WIDTH - 1 : 0] addr1,
        input wire [ADDR_WIDTH - 1 : 0] addr2,
        input wire wr_en1,
        input wire wr_en2,
        input wire [(1 << DATA_WIDTH) - 1 : 0] wr_data1,
        input wire [(1 << DATA_WIDTH) - 1 : 0] wr_data2,
        output wire [(1 << DATA_WIDTH) - 1 : 0] rd_data1,
        output wire [(1 << DATA_WIDTH) - 1 : 0] rd_data2
    );
        reg [(1 << DATA_WIDTH) - 1 : 0] mem [(1 << ADDR_WIDTH) - 1 : 0];
        reg [(1 << DATA_WIDTH) - 1 : 0] rd_data_reg1;
        reg [(1 << DATA_WIDTH) - 1 : 0] rd_data_reg2;
        assign rd_data1 = rd_data_reg1;
        assign rd_data2 = rd_data_reg2;
        always @(posedge clk) begin
            if(wr_en1) begin
                mem[addr1] <= wr_data1;
                rd_data_reg1 <= wr_data1;
            end else begin 
                rd_data_reg1 <= mem[addr1];
            end
        end
        always @(posedge clk) begin
            if(wr_en2) begin
                mem[addr2] <= wr_data2;
                rd_data_reg2 <= wr_data2;
            end else begin 
                rd_data_reg2 <= mem[addr2];
            end
        end
    endmodule
    module ram_t # (
        parameter DATA_WIDTH = 7,
        parameter ADDR_WIDTH = 10,
        parameter PARTITION_WIDTH = 4
    ) (
        input wire clk,
        input wire [ADDR_WIDTH - 1 : 0] addr1,
        input wire [ADDR_WIDTH - 1 : 0] addr2,
        input wire [ADDR_WIDTH - 1 : 0] offset_x1,
        input wire [ADDR_WIDTH - 1 : 0] offset_x2,
        input wire [ADDR_WIDTH - 1 : 0] offset_y1,
        input wire [ADDR_WIDTH - 1 : 0] offset_y2,
        input wire [(1 << PARTITION_WIDTH) - 1 : 0] wr_en1,
        input wire [(1 << PARTITION_WIDTH) - 1 : 0] wr_en2,
        input wire [(1 << DATA_WIDTH) - 1 : 0] wr_data1,
        input wire [(1 << DATA_WIDTH) - 1 : 0] wr_data2,
        output wire [(1 << DATA_WIDTH) - 1 : 0] rd_data1,
        output wire [(1 << DATA_WIDTH) - 1 : 0] rd_data2
    );
        reg [ADDR_WIDTH - 1 : 0] r_addr1;
        wire [ADDR_WIDTH - PARTITION_WIDTH - 1 : 0] p_addr1 [(1 << PARTITION_WIDTH) - 1 : 0];
        wire p_wr_en1 [(1 << PARTITION_WIDTH) - 1 : 0];
        wire [(1 << (DATA_WIDTH - PARTITION_WIDTH)) - 1 : 0] p_wr_data1 [(1 << PARTITION_WIDTH) - 1 : 0];
        wire [(1 << (DATA_WIDTH - PARTITION_WIDTH)) - 1 : 0] p_rd_data1 [(1 << PARTITION_WIDTH) - 1 : 0];
        wire [ADDR_WIDTH - PARTITION_WIDTH - 1 : 0] p_addr_next1, p_addr_curr1;
        wire [PARTITION_WIDTH - 1: 0] offset1;
        assign offset1 = r_addr1[PARTITION_WIDTH - 1 : 0]; 
        assign p_addr_next1 = &r_addr1[ADDR_WIDTH / 2 - 1 : PARTITION_WIDTH] ? {r_addr1[ADDR_WIDTH - 1 : ADDR_WIDTH / 2], {(ADDR_WIDTH / 2 - PARTITION_WIDTH){1'b0}}} : r_addr1[ADDR_WIDTH - 1 : PARTITION_WIDTH] + 1;
        assign p_addr_curr1 = r_addr1[ADDR_WIDTH - 1 : PARTITION_WIDTH];
        reg [ADDR_WIDTH - 1 : 0] r_addr2;
        wire [ADDR_WIDTH - PARTITION_WIDTH - 1 : 0] p_addr2 [(1 << PARTITION_WIDTH) - 1 : 0];
        wire p_wr_en2 [(1 << PARTITION_WIDTH) - 1 : 0];
        wire [(1 << (DATA_WIDTH - PARTITION_WIDTH)) - 1 : 0] p_wr_data2 [(1 << PARTITION_WIDTH) - 1 : 0];
        wire [(1 << (DATA_WIDTH - PARTITION_WIDTH)) - 1 : 0] p_rd_data2 [(1 << PARTITION_WIDTH) - 1 : 0];
        wire [ADDR_WIDTH - PARTITION_WIDTH - 1 : 0] p_addr_next2, p_addr_curr2;
        wire [PARTITION_WIDTH - 1: 0] offset2;
        assign offset2 = r_addr2[PARTITION_WIDTH - 1 : 0]; 
        assign p_addr_next2 = &r_addr2[ADDR_WIDTH / 2 - 1 : PARTITION_WIDTH] ? {r_addr2[ADDR_WIDTH - 1 : ADDR_WIDTH / 2], {(ADDR_WIDTH / 2 - PARTITION_WIDTH){1'b0}}} : r_addr2[ADDR_WIDTH - 1 : PARTITION_WIDTH] + 1;
        assign p_addr_curr2 = r_addr2[ADDR_WIDTH - 1 : PARTITION_WIDTH];
        always @(*) begin
            if((1 << (ADDR_WIDTH / 2)) - 1 - addr1[ADDR_WIDTH / 2 - 1 : 0] >= offset_x1) begin
                r_addr1[ADDR_WIDTH / 2 - 1 : 0] = addr1[ADDR_WIDTH / 2 - 1 : 0] + offset_x1;
            end else begin
                r_addr1[ADDR_WIDTH / 2 - 1 : 0] = offset_x1 - ((1 << (ADDR_WIDTH / 2)) - addr1[ADDR_WIDTH / 2 - 1 : 0]);
            end
            if((1 << (ADDR_WIDTH / 2)) - 1 - addr1[ADDR_WIDTH - 1 : ADDR_WIDTH / 2] >= offset_y1) begin
                r_addr1[ADDR_WIDTH - 1 : ADDR_WIDTH / 2] = addr1[ADDR_WIDTH - 1 : ADDR_WIDTH / 2] + offset_y1;
            end else begin
                r_addr1[ADDR_WIDTH - 1 : ADDR_WIDTH / 2] = offset_y1 - ((1 << (ADDR_WIDTH / 2)) - addr1[ADDR_WIDTH - 1 : ADDR_WIDTH / 2]);
            end
        end
        always @(*) begin
            if((1 << (ADDR_WIDTH / 2)) - 1 - addr2[ADDR_WIDTH / 2 - 1 : 0] >= offset_x2) begin
                r_addr2[ADDR_WIDTH / 2 - 1 : 0] = addr2[ADDR_WIDTH / 2 - 1 : 0] + offset_x2;
            end else begin
                r_addr2[ADDR_WIDTH / 2 - 1 : 0] = offset_x2 - ((1 << (ADDR_WIDTH / 2)) - addr2[ADDR_WIDTH / 2 - 1 : 0]);
            end
            if((1 << (ADDR_WIDTH / 2)) - 1 - addr2[ADDR_WIDTH - 1 : ADDR_WIDTH / 2] >= offset_y2) begin
                r_addr2[ADDR_WIDTH - 1 : ADDR_WIDTH / 2] = addr2[ADDR_WIDTH - 1 : ADDR_WIDTH / 2] + offset_y2;
            end else begin
                r_addr2[ADDR_WIDTH - 1 : ADDR_WIDTH / 2] = offset_y2 - ((1 << (ADDR_WIDTH / 2)) - addr2[ADDR_WIDTH - 1 : ADDR_WIDTH / 2]);
            end
        end
        genvar i;
        generate
            for(i = 0 ; i < (1 << PARTITION_WIDTH) ; i = i + 1) begin: gen_p_addr1
                assign p_addr1[i] = (i < offset1) ? p_addr_next1 : p_addr_curr1;
            end
            for(i = 0 ; i < (1 << PARTITION_WIDTH) ; i = i + 1) begin: gen_p_addr2
                assign p_addr2[i] = (i < offset2) ? p_addr_next2 : p_addr_curr2;
            end
            for(i = 0 ; i < (1 << PARTITION_WIDTH) ; i = i + 1) begin: gen_p_wr_wn1
                assign p_wr_en1[i] = wr_en1[(i < offset1) ?
                                            (i + (1 << PARTITION_WIDTH) - offset1) :
                                            (i - offset1)];
            end
            for(i = 0 ; i < (1 << PARTITION_WIDTH) ; i = i + 1) begin: gen_wr_en2
                assign p_wr_en2[i] = wr_en2[(i < offset2) ?
                                            (i + (1 << PARTITION_WIDTH) - offset2) :
                                            (i - offset2)];
            end
            for(i = 0 ; i < (1 << PARTITION_WIDTH) ; i = i + 1) begin: gen_p_wr_data1
                assign p_wr_data1[i] = wr_data1[((i < offset1) ? 
                                                (i + (1 << PARTITION_WIDTH) - offset1) : 
                                                (i - offset1)) << (DATA_WIDTH - PARTITION_WIDTH) +: 1 << (DATA_WIDTH - PARTITION_WIDTH)];
            end
            for(i = 0 ; i < (1 << PARTITION_WIDTH) ; i = i + 1) begin: gen_p_wr_data2
                assign p_wr_data2[i] = wr_data2[((i < offset2) ? 
                                                (i + (1 << PARTITION_WIDTH) - offset2) : 
                                                (i - offset2)) << (DATA_WIDTH - PARTITION_WIDTH) +: 1 << (DATA_WIDTH - PARTITION_WIDTH)];
            end
            for(i = 0 ; i < (1 << PARTITION_WIDTH) ; i = i + 1) begin: gen_ram
                p_ram_t # (.DATA_WIDTH((DATA_WIDTH - PARTITION_WIDTH)), .ADDR_WIDTH(ADDR_WIDTH - PARTITION_WIDTH)) ram (
                    .clk(clk),
                    .addr1(p_addr1[i]),
                    .addr2(p_addr2[i]),
                    .wr_en1(p_wr_en1[i]),
                    .wr_en2(p_wr_en2[i]),
                    .wr_data1(p_wr_data1[i]),
                    .wr_data2(p_wr_data2[i]),
                    .rd_data1(p_rd_data1[i]),
                    .rd_data2(p_rd_data2[i])
                );
            end
            for(i = 0 ; i < (1 << PARTITION_WIDTH) ; i = i + 1) begin: gen_p_rd_data1
                assign rd_data1[i << (DATA_WIDTH - PARTITION_WIDTH) +: 1 << (DATA_WIDTH - PARTITION_WIDTH)] = 
                    p_rd_data1[ (i < ((1 << (PARTITION_WIDTH)) - offset1)) ? 
                                (i + offset1) : 
                                (i - (1 << PARTITION_WIDTH) + offset1)];
            end
            for(i = 0 ; i < (1 << PARTITION_WIDTH) ; i = i + 1) begin: gen_p_rd_data2
                assign rd_data2[i << (DATA_WIDTH - PARTITION_WIDTH) +: 1 << (DATA_WIDTH - PARTITION_WIDTH)] = 
                    p_rd_data2[ (i < ((1 << (PARTITION_WIDTH)) - offset2)) ? 
                                (i + offset2) : 
                                (i - (1 << PARTITION_WIDTH) + offset2)];
            end
        endgenerate
    endmodule
	module data_provider_v1_0_S00_AXI #
	(
		// Users to add parameters here

		// User parameters ends
		// Do not modify the parameters beyond this line

		// Width of S_AXI data bus
		parameter integer C_S_AXI_DATA_WIDTH	= 32,
		// Width of S_AXI address bus
		parameter integer C_S_AXI_ADDR_WIDTH	= 6
	)
	(
		// Users to add ports here

		// User ports ends
		// Do not modify the ports beyond this line

		// Global Clock Signal
		input wire  S_AXI_ACLK,
		// Global Reset Signal. This Signal is Active LOW
		input wire  S_AXI_ARESETN,
		// Write address (issued by master, acceped by Slave)
		input wire [C_S_AXI_ADDR_WIDTH-1 : 0] S_AXI_AWADDR,
		// Write channel Protection type. This signal indicates the
    		// privilege and security level of the transaction, and whether
    		// the transaction is a data access or an instruction access.
		input wire [2 : 0] S_AXI_AWPROT,
		// Write address valid. This signal indicates that the master signaling
    		// valid write address and control information.
		input wire  S_AXI_AWVALID,
		// Write address ready. This signal indicates that the slave is ready
    		// to accept an address and associated control signals.
		output wire  S_AXI_AWREADY,
		// Write data (issued by master, acceped by Slave) 
		input wire [C_S_AXI_DATA_WIDTH-1 : 0] S_AXI_WDATA,
		// Write strobes. This signal indicates which byte lanes hold
    		// valid data. There is one write strobe bit for each eight
    		// bits of the write data bus.    
		input wire [(C_S_AXI_DATA_WIDTH/8)-1 : 0] S_AXI_WSTRB,
		// Write valid. This signal indicates that valid write
    		// data and strobes are available.
		input wire  S_AXI_WVALID,
		// Write ready. This signal indicates that the slave
    		// can accept the write data.
		output wire  S_AXI_WREADY,
		// Write response. This signal indicates the status
    		// of the write transaction.
		output wire [1 : 0] S_AXI_BRESP,
		// Write response valid. This signal indicates that the channel
    		// is signaling a valid write response.
		output wire  S_AXI_BVALID,
		// Response ready. This signal indicates that the master
    		// can accept a write response.
		input wire  S_AXI_BREADY,
		// Read address (issued by master, acceped by Slave)
		input wire [C_S_AXI_ADDR_WIDTH-1 : 0] S_AXI_ARADDR,
		// Protection type. This signal indicates the privilege
    		// and security level of the transaction, and whether the
    		// transaction is a data access or an instruction access.
		input wire [2 : 0] S_AXI_ARPROT,
		// Read address valid. This signal indicates that the channel
    		// is signaling valid read address and control information.
		input wire  S_AXI_ARVALID,
		// Read address ready. This signal indicates that the slave is
    		// ready to accept an address and associated control signals.
		output wire  S_AXI_ARREADY,
		// Read data (issued by slave)
		output wire [C_S_AXI_DATA_WIDTH-1 : 0] S_AXI_RDATA,
		// Read response. This signal indicates the status of the
    		// read transfer.
		output wire [1 : 0] S_AXI_RRESP,
		// Read valid. This signal indicates that the channel is
    		// signaling the required read data.
		output wire  S_AXI_RVALID,
		// Read ready. This signal indicates that the master can
    		// accept the read data and response information.
		input wire  S_AXI_RREADY
	);

	// AXI4LITE signals
	reg [C_S_AXI_ADDR_WIDTH-1 : 0] 	axi_awaddr;
	reg  	axi_awready;
	reg  	axi_wready;
	reg [1 : 0] 	axi_bresp;
	reg  	axi_bvalid;
	reg [C_S_AXI_ADDR_WIDTH-1 : 0] 	axi_araddr;
	reg  	axi_arready;
	reg [C_S_AXI_DATA_WIDTH-1 : 0] 	axi_rdata;
	reg [1 : 0] 	axi_rresp;
	reg  	axi_rvalid;

	// Example-specific design signals
	// local parameter for addressing 32 bit / 64 bit C_S_AXI_DATA_WIDTH
	// ADDR_LSB is used for addressing 32/64 bit registers/memories
	// ADDR_LSB = 2 for 32 bits (n downto 2)
	// ADDR_LSB = 3 for 64 bits (n downto 3)
	localparam integer ADDR_LSB = (C_S_AXI_DATA_WIDTH/32) + 1;
	localparam integer OPT_MEM_ADDR_BITS = 3;
	//----------------------------------------------
	//-- Signals for user logic register space example
	//------------------------------------------------
	//-- Number of Slave Registers 16
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg0;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg1;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg2;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg3;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg4;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg5;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg6;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg7;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg8;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg9;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg10;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg11;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg12;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg13;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg14;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg15;
	wire	 slv_reg_rden;
	wire	 slv_reg_wren;
	reg [C_S_AXI_DATA_WIDTH-1:0]	 reg_data_out;
	integer	 byte_index;

	// I/O Connections assignments

	assign S_AXI_AWREADY	= axi_awready;
	assign S_AXI_WREADY	= axi_wready;
	assign S_AXI_BRESP	= axi_bresp;
	assign S_AXI_BVALID	= axi_bvalid;
	assign S_AXI_ARREADY	= axi_arready;
	assign S_AXI_RDATA	= axi_rdata;
	assign S_AXI_RRESP	= axi_rresp;
	assign S_AXI_RVALID	= axi_rvalid;
	// Implement axi_awready generation
	// axi_awready is asserted for one S_AXI_ACLK clock cycle when both
	// S_AXI_AWVALID and S_AXI_WVALID are asserted. axi_awready is
	// de-asserted when reset is low.
	
	always @( posedge S_AXI_ACLK )
	begin
	  if ( S_AXI_ARESETN == 1'b0 )
	    begin
	      axi_awready <= 1'b0;
	    end 
	  else
	    begin    
	      if (~axi_awready && S_AXI_AWVALID && S_AXI_WVALID)
	        begin
	          // slave is ready to accept write address when 
	          // there is a valid write address and write data
	          // on the write address and data bus. This design 
	          // expects no outstanding transactions. 
	          axi_awready <= 1'b1;
	        end
	      else           
	        begin
	          axi_awready <= 1'b0;
	        end
	    end 
	end       

	// Implement axi_awaddr latching
	// This process is used to latch the address when both 
	// S_AXI_AWVALID and S_AXI_WVALID are valid. 

	always @( posedge S_AXI_ACLK )
	begin
	  if ( S_AXI_ARESETN == 1'b0 )
	    begin
	      axi_awaddr <= 0;
	    end 
	  else
	    begin    
	      if (~axi_awready && S_AXI_AWVALID && S_AXI_WVALID)
	        begin
	          // Write Address latching 
	          axi_awaddr <= S_AXI_AWADDR;
	        end
	    end 
	end       

	// Implement axi_wready generation
	// axi_wready is asserted for one S_AXI_ACLK clock cycle when both
	// S_AXI_AWVALID and S_AXI_WVALID are asserted. axi_wready is 
	// de-asserted when reset is low. 

	always @( posedge S_AXI_ACLK )
	begin
	  if ( S_AXI_ARESETN == 1'b0 )
	    begin
	      axi_wready <= 1'b0;
	    end 
	  else
	    begin    
	      if (~axi_wready && S_AXI_WVALID && S_AXI_AWVALID)
	        begin
	          // slave is ready to accept write data when 
	          // there is a valid write address and write data
	          // on the write address and data bus. This design 
	          // expects no outstanding transactions. 
	          axi_wready <= 1'b1;
	        end
	      else
	        begin
	          axi_wready <= 1'b0;
	        end
	    end 
	end       

	// Implement memory mapped register select and write logic generation
	// The write data is accepted and written to memory mapped registers when
	// axi_awready, S_AXI_WVALID, axi_wready and S_AXI_WVALID are asserted. Write strobes are used to
	// select byte enables of slave registers while writing.
	// These registers are cleared when reset (active low) is applied.
	// Slave register write enable is asserted when valid address and data are available
	// and the slave is ready to accept the write address and write data.
	wire [(1 << 8) - 1 : 0] rd_data;
    ram_t #(
        .ADDR_WIDTH(12),
        .DATA_WIDTH(8),
        .PARTITION_WIDTH(5)
    ) ram (
        .clk(S_AXI_ACLK),
        .addr1(slv_reg0[12 - 1 : 0]),
        .wr_en1({28'b0, {4{|slv_reg1}}}),
        .offset_x1(slv_reg2[12 - 1 : 0]),
        .offset_y1(slv_reg3[12 - 1 : 0]),
        .wr_data1({224'b0, slv_reg4}),
        .rd_data1(rd_data)
    );
	assign slv_reg_wren = axi_wready && S_AXI_WVALID && axi_awready && S_AXI_AWVALID;

	always @( posedge S_AXI_ACLK )
	begin
	  if ( S_AXI_ARESETN == 1'b0 )
	    begin
	      slv_reg0 <= 0;
	      slv_reg1 <= 0;
	      slv_reg2 <= 0;
	      slv_reg3 <= 0;
	      slv_reg4 <= 0;
	      slv_reg5 <= 0;
	      slv_reg6 <= 0;
	      slv_reg7 <= 0;
	      slv_reg8 <= 0;
	      slv_reg9 <= 0;
	      slv_reg10 <= 0;
	      slv_reg11 <= 0;
	      slv_reg12 <= 0;
	      slv_reg13 <= 0;
	      slv_reg14 <= 0;
	      slv_reg15 <= 0;
	    end 
	  else begin
	    if (slv_reg_wren)
	      begin
	        case ( axi_awaddr[ADDR_LSB+OPT_MEM_ADDR_BITS:ADDR_LSB] )
	          4'h0:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 0
	                slv_reg0[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	          4'h1:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 1
	                slv_reg1[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	          4'h2:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 2
	                slv_reg2[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	          4'h3:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 3
	                slv_reg3[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	          4'h4:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 4
	                slv_reg4[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	          4'h5:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 5
	                slv_reg5[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	          4'h6:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 6
	                slv_reg6[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	          4'h7:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 7
	                slv_reg7[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	          4'h8:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 8
	                slv_reg8[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	          4'h9:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 9
	                slv_reg9[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	          4'hA:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 10
	                slv_reg10[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	          4'hB:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 11
	                slv_reg11[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	          4'hC:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 12
	                slv_reg12[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	          4'hD:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 13
	                slv_reg13[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	          4'hE:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 14
	                slv_reg14[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	          4'hF:
	            for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
	              if ( S_AXI_WSTRB[byte_index] == 1 ) begin
	                // Respective byte enables are asserted as per write strobes 
	                // Slave register 15
	                slv_reg15[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
	              end  
	          default : begin
	                      slv_reg0 <= slv_reg0;
	                      slv_reg1 <= slv_reg1;
	                      slv_reg2 <= slv_reg2;
	                      slv_reg3 <= slv_reg3;
	                      slv_reg4 <= slv_reg4;
	                      slv_reg5 <= slv_reg5;
	                      slv_reg6 <= slv_reg6;
	                      slv_reg7 <= slv_reg7;
	                      slv_reg8 <= slv_reg8;
	                      slv_reg9 <= slv_reg9;
	                      slv_reg10 <= slv_reg10;
	                      slv_reg11 <= slv_reg11;
	                      slv_reg12 <= slv_reg12;
	                      slv_reg13 <= slv_reg13;
	                      slv_reg14 <= slv_reg14;
	                      slv_reg15 <= slv_reg15;
	                    end
	        endcase
	      end else begin
	      slv_reg0 <= slv_reg0;
                                    slv_reg1 <= slv_reg1;
                                    slv_reg2 <= slv_reg2;
                                    slv_reg3 <= slv_reg3;
                                    slv_reg4 <= slv_reg4;
                                    slv_reg5 <= rd_data[0 +: 32];
                                    slv_reg6 <= rd_data[32 +: 32];
                                    slv_reg7 <= rd_data[64 +: 32];
                                    slv_reg8 <= rd_data[96 +: 32];
                                    slv_reg9 <= rd_data[128 +: 32];
                                    slv_reg10 <= rd_data[160 +: 32];
                                    slv_reg11 <= rd_data[192 +: 32];
                                    slv_reg12 <= rd_data[224 +: 32];
                                    slv_reg13 <= slv_reg13;
                                    slv_reg14 <= slv_reg14;
                                    slv_reg15 <= slv_reg15;
	      end
	  end
	end    

	// Implement write response logic generation
	// The write response and response valid signals are asserted by the slave 
	// when axi_wready, S_AXI_WVALID, axi_wready and S_AXI_WVALID are asserted.  
	// This marks the acceptance of address and indicates the status of 
	// write transaction.

	always @( posedge S_AXI_ACLK )
	begin
	  if ( S_AXI_ARESETN == 1'b0 )
	    begin
	      axi_bvalid  <= 0;
	      axi_bresp   <= 2'b0;
	    end 
	  else
	    begin    
	      if (axi_awready && S_AXI_AWVALID && ~axi_bvalid && axi_wready && S_AXI_WVALID)
	        begin
	          // indicates a valid write response is available
	          axi_bvalid <= 1'b1;
	          axi_bresp  <= 2'b0; // 'OKAY' response 
	        end                   // work error responses in future
	      else
	        begin
	          if (S_AXI_BREADY && axi_bvalid) 
	            //check if bready is asserted while bvalid is high) 
	            //(there is a possibility that bready is always asserted high)   
	            begin
	              axi_bvalid <= 1'b0; 
	            end  
	        end
	    end
	end   

	// Implement axi_arready generation
	// axi_arready is asserted for one S_AXI_ACLK clock cycle when
	// S_AXI_ARVALID is asserted. axi_awready is 
	// de-asserted when reset (active low) is asserted. 
	// The read address is also latched when S_AXI_ARVALID is 
	// asserted. axi_araddr is reset to zero on reset assertion.

	always @( posedge S_AXI_ACLK )
	begin
	  if ( S_AXI_ARESETN == 1'b0 )
	    begin
	      axi_arready <= 1'b0;
	      axi_araddr  <= 32'b0;
	    end 
	  else
	    begin    
	      if (~axi_arready && S_AXI_ARVALID)
	        begin
	          // indicates that the slave has acceped the valid read address
	          axi_arready <= 1'b1;
	          // Read address latching
	          axi_araddr  <= S_AXI_ARADDR;
	        end
	      else
	        begin
	          axi_arready <= 1'b0;
	        end
	    end 
	end       

	// Implement axi_arvalid generation
	// axi_rvalid is asserted for one S_AXI_ACLK clock cycle when both 
	// S_AXI_ARVALID and axi_arready are asserted. The slave registers 
	// data are available on the axi_rdata bus at this instance. The 
	// assertion of axi_rvalid marks the validity of read data on the 
	// bus and axi_rresp indicates the status of read transaction.axi_rvalid 
	// is deasserted on reset (active low). axi_rresp and axi_rdata are 
	// cleared to zero on reset (active low).  
	always @( posedge S_AXI_ACLK )
	begin
	  if ( S_AXI_ARESETN == 1'b0 )
	    begin
	      axi_rvalid <= 0;
	      axi_rresp  <= 0;
	    end 
	  else
	    begin    
	      if (axi_arready && S_AXI_ARVALID && ~axi_rvalid)
	        begin
	          // Valid read data is available at the read data bus
	          axi_rvalid <= 1'b1;
	          axi_rresp  <= 2'b0; // 'OKAY' response
	        end   
	      else if (axi_rvalid && S_AXI_RREADY)
	        begin
	          // Read data is accepted by the master
	          axi_rvalid <= 1'b0;
	        end                
	    end
	end    

	// Implement memory mapped register select and read logic generation
	// Slave register read enable is asserted when valid address is available
	// and the slave is ready to accept the read address.
	assign slv_reg_rden = axi_arready & S_AXI_ARVALID & ~axi_rvalid;
	always @(*)
	begin
	      // Address decoding for reading registers
	      case ( axi_araddr[ADDR_LSB+OPT_MEM_ADDR_BITS:ADDR_LSB] )
	        4'h0   : reg_data_out <= slv_reg0;
	        4'h1   : reg_data_out <= slv_reg1;
	        4'h2   : reg_data_out <= slv_reg2;
	        4'h3   : reg_data_out <= slv_reg3;
	        4'h4   : reg_data_out <= slv_reg4;
	        4'h5   : reg_data_out <= slv_reg5;
	        4'h6   : reg_data_out <= slv_reg6;
	        4'h7   : reg_data_out <= slv_reg7;
	        4'h8   : reg_data_out <= slv_reg8;
	        4'h9   : reg_data_out <= slv_reg9;
	        4'hA   : reg_data_out <= slv_reg10;
	        4'hB   : reg_data_out <= slv_reg11;
	        4'hC   : reg_data_out <= slv_reg12;
	        4'hD   : reg_data_out <= slv_reg13;
	        4'hE   : reg_data_out <= slv_reg14;
	        4'hF   : reg_data_out <= slv_reg15;
	        default : reg_data_out <= 0;
	      endcase
	end

	// Output register or memory read data
	always @( posedge S_AXI_ACLK )
	begin
	  if ( S_AXI_ARESETN == 1'b0 )
	    begin
	      axi_rdata  <= 0;
	    end 
	  else
	    begin    
	      // When there is a valid read address (S_AXI_ARVALID) with 
	      // acceptance of read address by the slave (axi_arready), 
	      // output the read dada 
	      if (slv_reg_rden)
	        begin
	          axi_rdata <= reg_data_out;     // register read data
	        end   
	    end
	end    

	// Add user logic here

	// User logic ends

	endmodule
